library verilog;
use verilog.vl_types.all;
entity project01_test is
end project01_test;
