module ASmallerThanB(Z, Y, M);
	input Y, M;
	output Z;
	
	nor g(Z, Y, M);

endmodule
