library verilog;
use verilog.vl_types.all;
entity AGreaterThanB is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end AGreaterThanB;
